*TB
*-----------------------------------------------------------------
* HEAD
*-----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNWSW_CM_lpe.spi
#else
.include ../../../work/xsch/JNWSW_CM.spice
#endif
.option TNOM=27 GMIN=1e-15 reltol=1e-3 method=gear
.param TRF = 10p
.param AVDD = {vdda}
.param PERIOD_CLK = 1u
.param PW_CLK = PERIOD_CLK/2

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc {AVDD}
VCLK clk 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
VRESET reset 0 dc {AVDD} pwl 0 {AVDD} {PW_CLK*2} {AVDD} {PW_CLK*2 + 1n} 0
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names
VB0 b.0 b<0> dc 0
VB1 b.1 b<1> dc 0
VB2 b.2 b<2> dc 0
VB3 b.3 b<3> dc 0
VB4 b.4 b<4> dc 0

*- Bias current
IBPS 0 ibp dc 100n

* RC filter to calm the IDAC output
CDL IBN_DAC 0 10p
R1 IBN_DAC IBN_FILT 1k
VDAC IBN_FILT 0 dc 0.9

* The other bias currents
VI0 IBN_0 0 dc 0.9
VI1 IBN_1 0 dc 0.9
VI2 IBN_2 0 dc 0.9

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.save all
.save v(clk)
.save v(IBN_DAC)
.save v(IBN_FILT)
.save i(VDAC)
.save i(VI0)
.save i(VI1)
.save i(VI2)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

set fend = .raw

tran 125n 32u

write

quit


.endc

.end
